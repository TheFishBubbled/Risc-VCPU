module SingleCycleCPU(
        input CLK,                //????
        input Reset,              //????
        input reg[6:0] op,     
        input reg[2:0] funct3,  
        input reg[6:0] funct7,
        input reg[4:0] rs1,     
        input reg[4:0] rs2,     
        input reg[4:0] rd,     
        input reg[24:0] imm,    
        input reg [31:0] instr,  
        output [31:0] curPC      //????
    );


    wire [31:0] extend;    //???
  
   
    wire [31:0] DataOut;   //??????
    wire [1:0] cmp;      //?????
    //????
    wire PCSrc;
    wire [2:0] AluOp;
    wire AluSrc1;
    wire AluSrc2;
    wire RegWr;
    wire [1:0]RegDst;
    wire [2:0] ExtSel;
    wire Sign;
    wire [1:0] Digit;
    wire DataWr;
    wire immres;
    wire [31:0] AluOutput;
    wire[31:0] nextPC;
    wire[31:0]ReadData1;
    wire[31:0]ReadData2;
    wire[31:0]DB;

    PC pc(
        .CLK(CLK),       //??
        .Reset(Reset),   //??????
        .PCSrc(PCSrc),   //???????
        .AluOutput(AluOutput), //ALU????
        .curPC(curPC),    //???????
        .nextPC(nextPC)   //???
    );

    ControlUnit control(
        .cmp(cmp),        //?????
        .op(op),          //???
        .funct3(funct3),  //3????
        .funct7(funct7),  //7????
        .PCSrc(PCSrc),    //PC???????
        .AluOp(AluOp),    //ALU??
        .Alu1Src(AluSrc1),   //ALU1?
        .Alu2Src(AluSrc2),   //ALU2?
        .RegDst(RegDst),  //Rd??
        .RegWr(RegWr),    //Rd???
        .ExtSel(ExtSel),  //??????
        .Sign(Sign),      //???????
        .Digit(Digit),    //????
        .DataWr(DataWr),  //??????
        .immres(immres)   //rd????imm??????
    );

    ALU alu(
        .ALUSrc1(AluSrc1),     //???1??
        .ALUSrc2(AluSrc2),     //???2??
        .ReadData1(ReadData1), //rs1???????
        .ReadData2(ReadData2), //rs2???????
        .extend(extend),       //??????
        .PC(curPC),            //????????????
        .AluOp(AluOp),         //ALU???
        .cmp(cmp),             //???????
        .AluOutput(AluOutput),  //ALU????
	.Sign(Sign)
    );
/*
    InsMEM insmem(
        .curPC(curPC),   //PC?
        .op(op),         //?????
        .funct3(funct3), //3??????
        .funct7(funct7), //7??????
        .rs1(rs1),       //rs2????
        .rs2(rs2),       //rs2????
        .rd(rd),         //rd????
        .imm(imm),       //???????extend??????
        .instr(instr)    //????32???
    );
*/

    Extend ext(
        .imm(imm),        //?????
        .ExtSel(ExtSel),  //????
        .extend(extend)   //??????
    );

    RegisterFile regfile(
        .CLK(CLK),         //??
        .immres(immres),   //?????????
        .rs1(rs1),         //rs1?????????
        .rs2(rs2),         //rs2?????????
        .WriteReg(rd),
        .AluOutput(AluOutput), //ALU??
        .extend(extend),       //imm?????
        .Datain(DataOut),      //?????
        .PC(curPC),            //??PC?
        .cmp(cmp),             //?????
        .RegDst(RegDst),       //????????
        .RegWr(RegWr),         //???????1??????????
        .DB(DB),               //??????
        .ReadData1(ReadData1), //rs1?????????
        .ReadData2(ReadData2)  //rs2?????????
    );

    DataMEM datamem(
        .DataWr(DataWr), //??????
        .Digit(Digit), //?????00?8??01?16??10?32?
        .CLK(CLK),     //?????????
        .DAddr(AluOutput),  //????
        .DataIn(ReadData2), //????
        .DataOut(DataOut), //????
	.pc(curPC)
    );

endmodule